.title KiCad schematic
J2 Net-_J2-Pad1_ Net-_J1-Pad1_ Net-_J2-Pad3_ Conn_01x03
J3 Net-_J2-Pad1_ Net-_J2-Pad3_ Net-_J1-Pad2_ Net-_J1-Pad3_ Net-_J1-Pad4_ NC_01 Net-_J1-Pad6_ Net-_J1-Pad5_ Net-_J1-Pad7_ Net-_J1-Pad8_ Conn_02x05_Odd_Even
J1 Net-_J1-Pad1_ Net-_J1-Pad2_ Net-_J1-Pad3_ Net-_J1-Pad4_ Net-_J1-Pad5_ Net-_J1-Pad6_ Net-_J1-Pad7_ Net-_J1-Pad8_ RJ45
.end
